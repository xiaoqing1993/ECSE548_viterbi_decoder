*** SPICE deck for cell inv_1x{sch} from library Project
*** Created on Wed Oct 11, 2006 19:45:21
*** Last revised on Mon Mar 12, 2007 05:28:50
*** Written on Thu Dec 01, 2016 02:41:27 by Electric VLSI Design System, 
*version 8.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
.OPTIONS NOMOD NOPAGE
*CMOS/BULK-NWELL (PRELIMINARY PARAMETERS)
.OPTIONS NOMOD DEFL=3UM DEFW=3UM DEFAD=70P DEFAS=70P LIMPTS=1000
+ITL5=0 RELTOL=0.01 ABSTOL=500PA VNTOL=500UV LVLTIM=2
+LVLCOD=1
.MODEL N NMOS LEVEL=1
+KP=60E-6 VTO=0.7 GAMMA=0.3 LAMBDA=0.05 PHI=0.6
+LD=0.4E-6 TOX=40E-9 CGSO=2.0E-10 CGDO=2.0E-10 CJ=.2MF/M^2
.MODEL P PMOS LEVEL=1
+KP=20E-6 VTO=0.7 GAMMA=0.4 LAMBDA=0.05 PHI=0.6
+LD=0.6E-6 TOX=40E-9 CGSO=3.0E-10 CGDO=3.0E-10 CJ=.2MF/M^2
.MODEL DIFFCAP D CJO=.2MF/M^2

.global gnd vdd

*** TOP LEVEL CELL: inv_1x{sch}
Mnmos@0 y a gnd gnd N L=0.6U W=2.1U
Mpmos@0 vdd a y vdd P L=0.6U W=3U
.END
