*** SPICE deck for cell adder6_ksa{sch} from library Project
*** Created on Thu Nov 24, 2016 15:28:06
*** Last revised on Sat Nov 26, 2016 03:05:07
*** Written on Thu Dec 01, 2016 02:38:54 by Electric VLSI Design System,
*version 8.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* DATE: Jan  7/09
* LOT: T89Y                  WAF: 7103
* Temperature_parameters=Default
.MODEL N NMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 1.41E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = 0.6490078
+K1      = 0.8791883      K2      = -0.0987192     K3      = 30.3743151
+K3B     = -8.9028418     W0      = 1E-8           NLX     = 1E-9
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.7760383      DVT1    = 0.3617427      DVT2    = -0.4947423
+U0      = 448.0056882    UA      = 1E-13          UB      = 1.232756E-18
+UC      = 1.919293E-12   VSAT    = 1.853447E5     A0      = 0.6608042
+AGS     = 0.1481249      B0      = 2.156839E-6    B1      = 5E-6
+KETA    = -5.124492E-3   A1      = 2.16677E-6     A2      = 0.3
+RDSW    = 1.221635E3     PRWG    = 0.1064777      PRWB    = 0.0440597
+WR      = 1              WINT    = 2.288199E-7    LINT    = 9.639076E-8
+XL      = 1E-7           XW      = 0              DWG     = -1.520128E-9
+DWB     = 4.808525E-8    VOFF    = 0              NFACTOR = 1.230707
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 7.012161E-3    ETAB    = 4.092429E-4
+DSUB    = 0.2049812      PCLM    = 2.8412194      PDIBLC1 = 9.256485E-4
+PDIBLC2 = 2.355065E-3    PDIBLCB = -2.620257E-3   DROUT   = 0.0454337
+PSCBE1  = 6.464275E8     PSCBE2  = 2.427079E-4    PVAG    = 0
+DELTA   = 0.01           RSH     = 87.7           MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 1.79E-10       CGSO    = 1.79E-10       CGBO    = 1E-9
+CJ      = 4.136412E-4    PB      = 0.8475328      MJ      = 0.4294826
+CJSW    = 3.231457E-10   PBSW    = 0.8            MJSW    = 0.1846141
+CJSWG   = 1.64E-10       PBSWG   = 0.8            MJSWG   = 0.1846141
+CF      = 0              PVTH0   = -0.0466277     PRDSW   = 500
+PK2     = -0.0737963     WKETA   = -0.0147458     LKETA   = -2.029778E-3    )
*
.MODEL P PMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 1.41E-8
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = -0.9152268
+K1      = 0.553472       K2      = 7.871921E-3    K3      = 22.5354609
+K3B     = -1.1112458     W0      = 2.03458E-6     NLX     = 1.722913E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 1.2139827      DVT1    = 0.3310703      DVT2    = -0.0693525
+U0      = 201.3603195    UA      = 2.408572E-9    UB      = 1E-21
+UC      = -1E-10         VSAT    = 8.995975E4     A0      = 0.8936587
+AGS     = 0.0900735      B0      = 7.860659E-8    B1      = 3.278183E-9
+KETA    = -4.865785E-3   A1      = 2.887338E-4    A2      = 0.6177492
+RDSW    = 3E3            PRWG    = -0.0301252     PRWB    = -0.0443005
+WR      = 1              WINT    = 2.76783E-7     LINT    = 1.184609E-7
+XL      = 1E-7           XW      = 0              DWG     = 6.999518E-10
+DWB     = -8.293887E-9   VOFF    = -0.0727048     NFACTOR = 1.0504728
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 3.502584E-4    ETAB    = -0.2
+DSUB    = 1              PCLM    = 2.3553185      PDIBLC1 = 0.0614112
+PDIBLC2 = 2.759101E-3    PDIBLCB = -0.0320372     DROUT   = 0.2875724
+PSCBE1  = 1E8            PSCBE2  = 3.337278E-9    PVAG    = 9.077394E-4
+DELTA   = 0.01           RSH     = 110.4          MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 2.1E-10        CGSO    = 2.1E-10        CGBO    = 1E-9
+CJ      = 7.174866E-4    PB      = 0.9112434      MJ      = 0.4943334
+CJSW    = 2.179589E-10   PBSW    = 0.99           MJSW    = 0.2586376
+CJSWG   = 6.4E-11        PBSWG   = 0.99           MJSWG   = 0.2586376
+CF      = 0              PVTH0   = 5.98016E-3     PRDSW   = 14.8598424
+PK2     = 3.73981E-3     WKETA   = 0.0119588      LKETA   = -0.0101021      )
*

*** CELL: and3_1x{sch}
.SUBCKT and3_1x a b c y
Mnmos@0 net@9 b net@45 gnd N L=0.6U W=2.4U
Mnmos@1 net@1 c net@9 gnd N L=0.6U W=2.4U
Mnmos@3 y net@1 gnd gnd N L=0.6U W=2.1U
Mnmos@4 net@45 a gnd gnd N L=0.6U W=2.4U
Mpmos@0 vdd c net@1 vdd P L=0.6U W=1.8U
Mpmos@1 vdd net@1 y vdd P L=0.6U W=3U
Mpmos@2 vdd a net@1 vdd P L=0.6U W=1.8U
Mpmos@3 vdd b net@1 vdd P L=0.6U W=1.8U
.ENDS and3_1x

*** CELL: inv_1x{sch}
.SUBCKT inv_1x a y
Mnmos@0 y a gnd gnd N L=0.6U W=2.1U
Mpmos@0 vdd a y vdd P L=0.6U W=3U
.ENDS inv_1x

*** CELL: mux2_c_1x{sch}
.SUBCKT mux2_c_1x d0 d1 s y
Mnmos@0 net@3 d1 gnd gnd N L=0.6U W=1.8U
Mnmos@1 net@4 d0 gnd gnd N L=0.6U W=1.8U
Mnmos@2 net@5 s net@3 gnd N L=0.6U W=1.8U
Mnmos@3 net@5 sb net@4 gnd N L=0.6U W=1.8U
Mnmos@4 y net@5 gnd gnd N L=0.6U W=2.1U
Mnmos@5 sb s gnd gnd N L=0.6U W=1.8U
Mpmos@0 net@15 sb net@5 vdd P L=0.6U W=2.7U
Mpmos@1 vdd d1 net@15 vdd P L=0.6U W=2.7U
Mpmos@2 net@12 s net@5 vdd P L=0.6U W=2.7U
Mpmos@3 vdd d0 net@12 vdd P L=0.6U W=2.7U
Mpmos@4 vdd net@5 y vdd P L=0.6U W=3U
Mpmos@5 vdd s sb vdd P L=0.6U W=2.7U
.ENDS mux2_c_1x

*** CELL: mux6{sch}
.SUBCKT mux6 d0[0] d0[1] d0[2] d0[3] d0[4] d0[5] d1[0] d1[1] d1[2] d1[3]
+d1[4] d1[5] s y[0] y[1] y[2] y[3] y[4] y[5]
Xmux2_c_1@0 d0[0] d1[0] s y[0] mux2_c_1x
Xmux2_c_1@1 d0[1] d1[1] s y[1] mux2_c_1x
Xmux2_c_1@2 d0[2] d1[2] s y[2] mux2_c_1x
Xmux2_c_1@3 d0[3] d1[3] s y[3] mux2_c_1x
Xmux2_c_1@4 d0[4] d1[4] s y[4] mux2_c_1x
Xmux2_c_1@5 d0[5] d1[5] s y[5] mux2_c_1x
.ENDS mux6

*** CELL: and2_1x{sch}
.SUBCKT and2_1x a b y
Mnmos@0 net@2 b net@1 gnd N L=0.6U W=1.8U
Mnmos@1 net@1 a gnd gnd N L=0.6U W=1.8U
Mnmos@2 y net@2 gnd gnd N L=0.6U W=2.1U
Mpmos@0 vdd b net@2 vdd P L=0.6U W=1.8U
Mpmos@1 vdd a net@2 vdd P L=0.6U W=1.8U
Mpmos@2 vdd net@2 y vdd P L=0.6U W=3U
.ENDS and2_1x

*** CELL: xor2_1x{sch}
.SUBCKT xor2_1x a b y
Mnmos@0 net@3 a gnd gnd N L=0.6U W=4.2U
Mnmos@1 net@4 ab gnd gnd N L=0.6U W=4.2U
Mnmos@2 y b net@3 gnd N L=0.6U W=4.2U
Mnmos@3 y bb net@4 gnd N L=0.6U W=4.2U
Mnmos@4 bb b gnd gnd N L=0.6U W=1.8U
Mnmos@5 ab a gnd gnd N L=0.6U W=1.8U
Mpmos@0 net@7 b y vdd P L=0.6U W=6U
Mpmos@1 vdd ab net@7 vdd P L=0.6U W=6U
Mpmos@2 net@8 bb y vdd P L=0.6U W=6U
Mpmos@3 vdd a net@8 vdd P L=0.6U W=6U
Mpmos@4 vdd b bb vdd P L=0.6U W=2.7U
Mpmos@5 vdd a ab vdd P L=0.6U W=2.7U
.ENDS xor2_1x

*** CELL: bit_prop_gen{sch}
.SUBCKT bit_prop_gen A B G P
Xand2_1x@0 A B G and2_1x
Xxor2_1x@0 A B P xor2_1x
.ENDS bit_prop_gen

*** CELL: a2o1_1x{sch}
.SUBCKT a2o1_1x a b c y
Mnmos@0 net@19 a gnd gnd N L=0.6U W=1.8U
Mnmos@1 net@0 b net@19 gnd N L=0.6U W=1.8U
Mnmos@2 net@0 c gnd gnd N L=0.6U W=1.8U
Mnmos@3 y net@0 gnd gnd N L=0.6U W=2.1U
Mpmos@0 net@11 c net@0 vdd P L=0.6U W=2.7U
Mpmos@1 vdd b net@11 vdd P L=0.6U W=2.7U
Mpmos@2 vdd a net@11 vdd P L=0.6U W=2.7U
Mpmos@3 vdd net@0 y vdd P L=0.6U W=3U
.ENDS a2o1_1x

*** CELL: group_gen{sch}
.SUBCKT group_gen G0 G1 G2 P1
Xa2o1_1x@0 G0 P1 G1 G2 a2o1_1x
.ENDS group_gen

*** CELL: group_prop_gen{sch}
.SUBCKT group_prop_gen G0 G1 G2 P0 P1 P2
Xa2o1_1x@0 G0 P1 G1 G2 a2o1_1x
Xand2_1x@0 P0 P1 P2 and2_1x
.ENDS group_prop_gen

*** CELL: six_bit_kogge_stone_adder{sch}
.SUBCKT six_bit_kogge_stone_adder A[0] A[1] A[2] A[3] A[4] A[5] B[0] B[1]
+B[2] B[3] B[4] B[5] S[0] S[1] S[2] S[3] S[4] S[5]
Xbit_prop@0 A[0] B[0] net@0 P[0] bit_prop_gen
Xbit_prop@1 A[1] B[1] net@2 P[1] bit_prop_gen
Xbit_prop@2 A[2] B[2] net@4 P[2] bit_prop_gen
Xbit_prop@3 A[3] B[3] net@6 P[3] bit_prop_gen
Xbit_prop@4 A[4] B[4] net@144 P[4] bit_prop_gen
Xbit_prop@5 A[5] B[5] bit_prop@5_G P[5] bit_prop_gen
Xgroup_ge@0 gnd net@0 net@71 P[0] group_gen
Xgroup_ge@1 gnd net@20 net@143 net@21 group_gen
Xgroup_ge@2 net@71 net@18 net@120 net@19 group_gen
Xgroup_ge@3 gnd net@26 net@119 net@27 group_gen
Xgroup_ge@4 net@71 net@24 net@115 net@25 group_gen
Xgroup_pr@0 net@2 net@4 net@18 P[1] P[2] net@19 group_prop_gen
Xgroup_pr@1 net@0 net@2 net@20 P[0] P[1] net@21 group_prop_gen
Xgroup_pr@2 net@4 net@6 net@141 P[2] P[3] net@142 group_prop_gen
Xgroup_pr@3 net@6 net@144 net@14 P[3] P[4] net@15 group_prop_gen
Xgroup_pr@5 net@20 net@141 net@26 net@21 net@142 net@27 group_prop_gen
Xgroup_pr@6 net@18 net@14 net@24 net@19 net@15 net@25 group_prop_gen
Xxor2_1x@0 net@115 P[5] S[5] xor2_1x
Xxor2_1x@4 net@119 P[4] S[4] xor2_1x
Xxor2_1x@5 net@120 P[3] S[3] xor2_1x
Xxor2_1x@6 net@143 P[2] S[2] xor2_1x
Xxor2_1x@7 net@71 P[1] S[1] xor2_1x
Xxor2_1x@8 gnd P[0] S[0] xor2_1x
.ENDS six_bit_kogge_stone_adder

.global gnd vdd

*** TOP LEVEL CELL: adder6_ksa{sch}
Xand3_1x@0 b[5] net@21 a[5] net@19 and3_1x
Xand3_1x@1 net@22 s[5] net@24 net@20 and3_1x
Xinv_1x@0 s[5] net@21 inv_1x
Xinv_1x@1 a[5] net@24 inv_1x
Xinv_1x@2 b[5] net@22 inv_1x
Xmux6@0 s[0] s[1] s[2] s[3] s[4] s[5] gnd gnd gnd gnd gnd vdd net@19
+net@15[0] net@15[1] net@15[2] net@15[3] net@15[4] net@15[5] mux6
Xmux6@1 net@15[0] net@15[1] net@15[2] net@15[3] net@15[4] net@15[5] vdd vdd
+vdd vdd vdd gnd net@20 y[0] y[1] y[2] y[3] y[4] y[5] mux6
Xsix_bit_@0 a[0] a[1] a[2] a[3] a[4] a[5] b[0] b[1] b[2] b[3] b[4] b[5] s[0]
+s[1] s[2] s[3] s[4] s[5] six_bit_kogge_stone_adder

*** Load - KS avg
C1 y[5] 0 38.59F
C2 y[4] 0 38.59F
C3 y[3] 0 38.59F
C4 y[2] 0 38.59F
C5 y[1] 0 38.59F
C6 y[0] 0 38.59F

*** Test voltages
vdd VDD 0 DC 5
V1 a[0] 0 PULSE(0 5 100n 0.1n 0.1n 100n 200n 2056)
V2 a[1] 0 PULSE(0 5 200n 0.1n 0.1n 200n 400n 1024)
V3 a[2] 0 PULSE(0 5 400n 0.1n 0.1n 400n 800n 512)
V4 a[3] 0 PULSE(0 5 800n 0.1n 0.1n 800n 1600n 256)
V5 a[4] 0 PULSE(0 5 1600n 0.1n 0.1n 1600n 3200n 128)
V6 a[5] 0 PULSE(0 5 3200n 0.1n 0.1n 3200n 6400n 64)
V7 b[0] 0 PULSE(0 5 6400n 0.1n 0.1n 6400n 12800n 32)
V8 b[1] 0 PULSE(0 5 12800n 0.1n 0.1n 12800n 25600n 16)
V9 b[2] 0 PULSE(0 5 25600n 0.1n 0.1n 25600n 51200n 8)
V10 b[3] 0 PULSE(0 5 51200n 0.1n 0.1n 51200n 102400n 4)
V11 b[4] 0 PULSE(0 5 102400n 0.1n 0.1n 102400n 204800n 2)
V12 b[5] 0 PULSE(0 5 204800n 0.1n 0.1n 204800n 409600n 1)
.tran 409.6u
.END
