library verilog;
use verilog.vl_types.all;
entity six_bit_kogge_stone_adder_vlg_vec_tst is
end six_bit_kogge_stone_adder_vlg_vec_tst;
